library verilog;
use verilog.vl_types.all;
entity UAL_vlg_vec_tst is
end UAL_vlg_vec_tst;
